LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY T_TRIGGER IS 

PORT(
CLK, T: IN STD_LOGIC;
CLEAR: IN STD_LOGIC;
S1: INOUT STD_LOGIC;
S2: INOUT STD_LOGIC

);
END T_TRIGGER;


ARCHITECTURE BEHAVE OF T_TRIGGER IS 

BEGIN

 
PROCESS(CLK, CLEAR)
BEGIN

IF(S1 = 'U')THEN
	S1 <= '0';
	S2 <= '1';
END IF;

IF(CLEAR = '1')THEN
	S1 <= '0';
	S2 <= '1';

ELSIF(CLK'EVENT AND CLK = '1' AND T = '1')THEN

	S1 <= NOT(S1);
	S2 <= NOT(S2);
	
END IF;

END PROCESS;


END BEHAVE;