LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY myDFF IS

PORT(
CLK: IN STD_LOGIC;
D: INOUT STD_LOGIC;
ENABLE: IN STD_LOGIC;
OUTPUT: INOUT STD_LOGIC

);

END myDFF;



ARCHITECTURE BEHAVE OF myDFF IS 

BEGIN



PROCESS(CLK)BEGIN	

	IF(ENABLE = '1')THEN
		IF(clk'EVENT AND CLK = '1')THEN

			OUTPUT <= NOT(OUTPUT);

		END IF;

	END IF;

	IF(OUTPUT = 'U')THEN
		OUTPUT <= '0';

	END IF;

END PROCESS;

END BEHAVE;