LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

--
--	Pseudo random number generator - SAS
--


Entity RandomNumber is
port(

	requestLine: in std_logic;
	newData: out std_logic := '0';
	lastNumberGenerated: inout natural := 500;
	newNumberGenerated: inout natural := 500;
	dataLine: out std_logic_vector(11 downto 0);
	min: in std_logic_vector(11 downto 0);
	max: in std_logic_vector(11 downto 0)
	
);
End RandomNumber;


Architecture hardRN of RandomNumber is 

signal a: natural := 397204094;
signal m: natural := 1073741823;
signal c: natural := 0; 

--signal lastNumberGenerated: natural;
--signal newNumberGenerated: natural;

signal min_n : natural range 0 to 900;															--minimum number that can be generated by the algorithm
signal max_n: natural range 0 to 1440;															--maximimum number that can be generated by the algorithm

begin 

	--
	--	A new number will be generated when is requested over requestLine
	--
	min_n <= to_integer(unsigned(min));
	max_n <= to_integer(unsigned(max));
	
	new_number: process(requestLine)
		
		begin
		if(rising_edge(requestLine))then	
			
			newNumberGenerated <= integer(((lastNumberGenerated * a + c) mod m) mod max_n);
	
			lastNumberGenerated <= integer(newNumberGenerated * (max_n - min_n)/max_n) + min_n;
			
			dataLine <= std_logic_vector(to_unsigned( lastNumberGenerated, dataLine'length ));
			
			newData <= not(newData);

		end if;
	
	end process;
	
end hardRN;