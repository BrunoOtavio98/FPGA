LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARADOR IS 
GENERIC(N: INTEGER := 32);

PORT(

INPUT: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
CTE: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);

OUTPUT_EQUAL: OUT STD_LOGIC;
OUTPUT_GREATER: OUT STD_LOGIC

);
END COMPARADOR;

ARCHITECTURE BEHAVE OF COMPARADOR IS
BEGIN 
OUTPUT_EQUAL <= '1' WHEN (INPUT = CTE) ELSE
					 '0';
					 
OUTPUT_GREATER <= '1' WHEN (INPUT > CTE) ELSE
						 '0';
END BEHAVE;